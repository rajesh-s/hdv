package pack;
`include "env_adder_packet.sv"
`include "env_adder_generator.sv"
`include "env_adder_driver.sv"
`include "env_adder_intf.sv"
`include "env_adder_coverage.sv"// This inclusion is dependent on the position.
`include "env_adder.sv"
`include "env_adder_monitor.sv"
`include "env_adder_scoreboard.sv"
`include "env_adder_environment.sv"
`include "env_adder_test.sv"
endpackage
