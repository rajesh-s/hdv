module fourth;
struct
{
	integer payload;
	bit [11:0] data;
	shortint crc;
} fourth;
endmodule

