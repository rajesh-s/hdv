class base;
int j = 7;
task print();
begin
	$display("%d",j);
end
endtask
endclass
