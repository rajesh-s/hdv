module adder(input [15:0] a,b, output logic [16:0] sum);
assign sum = a + b;
endmodule
