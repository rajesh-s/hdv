module array;
bit [0:4][31:0] pack;
initial
	//pack[6] = 11;
	$display("array [] = %0d",pack[5]);
endmodule
