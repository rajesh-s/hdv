module rhs_lhs;
int a =9;
initial
begin
a= a;
$display("%d",a);
end
endmodule
