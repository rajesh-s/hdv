module race_condition;

initial 
  $display(" Initial 1");

initial 
  $display(" Initial 2");

initial 
  $display(" Initial 3");
endmodule
